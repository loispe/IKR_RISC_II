--
-- VHDL Architecture raro_ikr_risc_II_lib.man_clk_sim.behav
--
-- Created:
--          by - kntntply.meyer (pc091)
--          at - 14:37:48 07/13/22
--
-- using Mentor Graphics HDL Designer(TM) 2020.2 Built on 12 Apr 2020 at 11:28:22
--
ARCHITECTURE behav OF man_clk_sim IS
BEGIN
  sel_clk <= '0';
  man_clk <= '0';
END ARCHITECTURE behav;

