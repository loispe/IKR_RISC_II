--
-- VHDL Architecture raro_ikr_risc_II_lib.step_me.behav
--
-- Created:
--          by - lspetrck.meyer (pc091)
--          at - 14:17:51 05/25/22
--
-- using Mentor Graphics HDL Designer(TM) 2020.2 Built on 12 Apr 2020 at 11:28:22
--
ARCHITECTURE behav OF step_me IS
BEGIN
  rME_in <= rALU_out;
END ARCHITECTURE behav;

