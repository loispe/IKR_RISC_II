--
-- vhdl architecture raro_ikr_risc_ii_lib.man_clk_sim.behav
--
-- created:
--          by - kntntply.meyer (pc091)
--          at - 14:37:48 07/13/22
--
-- using mentor graphics hdl designer(tm) 2020.2 built on 12 apr 2020 at 11:28:22
--
architecture behav of man_clk_sim is
begin
  sel_clk <= '0';
  man_clk <= '0';
end architecture behav;

